module SEGMENT_ABS_ADD(CLK, A,B, N_Reset, SEG_COM, SEG_DATA);

input CLK, N_Reset;
input [3:0] A;
input [3:0] B;
output [7:0] SEG_COM, SEG_DATA;
wire [3:0] I;
wire C_OUT;
LAB03_4BIT_ABS H1(A,B,C_OUT,I);
wire [9:0] BCD_OUT; 
wire A1,B1,C1,D1,E1,F1,G1,A2,B2,C2,D2,E2,F2,G2;
//LAB04_BINTOBCD(B,P);
//LAB04_BCD_TO_7SEGMENT(BCD,A,B,C,D,E,F,G)
LAB04_BINTOBCD U1(I,BCD_OUT); 
LAB04_BCD_TO_7SEGMENT U2(BCD_OUT[3:0],A1,B1,C1,D1,E1,F1,G1);
LAB04_BCD_TO_7SEGMENT U3(BCD_OUT[7:4],A2,B2,C2,D2,E2,F2,G2);

LAB04_7SEG_CTRL U4(CLK, N_Reset, {A1,B1,C1,D1,E1,F1,G1},{A2,B2,C2,D2,E2,F2,G2}, 0,0,0,0,0,0,SEG_COM, SEG_DATA); 

endmodule