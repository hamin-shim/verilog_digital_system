

module LAB05_D_FF(CLK, D, Q, NQ);
  input CLK, D;
  output Q, NQ;
  wire w1, w2, w3, w4;
  LAB05_SR_LATCH L1(.S(w4), .R(CLK), .Q(w1), .NQ(w2));
  LAB05_SR_LATCH L2(.S(w2&CLK), .R(D), .Q(w3), .NQ(w4));
  LAB05_SR_LATCH L3(.S(w2), .R(w3), .Q(Q), .NQ(NQ));
endmodule
