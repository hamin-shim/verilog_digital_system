`timescale 10ns/1ps

module LAB03_HALFADDER_TB;

	reg A;
	reg B;

	
	LAB03_HALFADDER U1(A,B,Y,Z);
	initial begin
		A<=0;B<=0;
		#10 A<=0;B<=1;
		#10 A<=1;B<=0;
		#10 A<=1;B<=1;
	end
    
endmodule